library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is   
  port(
    clk     : in  std_logic;
    address : in  std_logic_vector(146 downto 0);
    data1   : out std_logic;
    data2   : out std_logic;
    data3   : out std_logic;
    data4   : out std_logic;
    data5   : out std_logic;
    data6   : out std_logic
  );       
end entity;

architecture RTL of rom is
  subtype byte is std_logic;
  type memory  is array (146 downto 0) of byte;

  constant vector1 : memory := 
  (
    0   =>'0', 1   =>'1', 2   =>'1', 3   =>'1', 4   =>'0', 5   =>'0', 6   =>'1', 7   =>'0', 8   =>'1', 9   =>'0', 
    10  =>'1', 11  =>'1', 12  =>'0', 13  =>'1', 14  =>'0', 15  =>'0', 16  =>'0', 17  =>'1', 18  =>'0', 19  =>'1', 
    20  =>'1', 21  =>'1', 22  =>'0', 23  =>'0', 24  =>'1', 25  =>'0', 26  =>'1', 27  =>'0', 28  =>'1', 29  =>'0', 
    30  =>'1', 31  =>'0', 32  =>'0', 33  =>'1', 34  =>'0', 35  =>'0', 36  =>'0', 37  =>'1', 38  =>'1', 39  =>'0', 
    40  =>'0', 41  =>'1', 42  =>'1', 43  =>'0', 44  =>'0', 45  =>'0', 46  =>'1', 47  =>'1', 48  =>'0', 49  =>'0',
    50  =>'1', 51  =>'1', 52  =>'0', 53  =>'0', 54  =>'1', 55  =>'1', 56  =>'1', 57  =>'0', 58  =>'1', 59  =>'0', 
    60  =>'0', 61  =>'1', 62  =>'0', 63  =>'1', 64  =>'1', 65  =>'1', 66  =>'0', 67  =>'0', 68  =>'1', 69  =>'1',
    70  =>'0', 71  =>'0', 72  =>'0', 73  =>'1', 74  =>'0', 75  =>'1', 76  =>'1', 77  =>'0', 78  =>'1', 79  =>'0', 
    80  =>'1', 81  =>'0', 82  =>'1', 83  =>'0', 84  =>'0', 85  =>'1', 86  =>'1', 87  =>'0', 88  =>'1', 89  =>'0',
    90  =>'1', 91  =>'0', 92  =>'1', 93  =>'1', 94  =>'0', 95  =>'1', 96  =>'1', 97  =>'1', 98  =>'0', 99  =>'0',
    100 =>'0', 101 =>'0', 102 =>'1', 103 =>'1', 104 =>'1', 105 =>'1', 106 =>'0', 107 =>'0', 108 =>'1', 109 =>'1', 
    110 =>'1', 111 =>'1', 112 =>'0', 113 =>'0', 114 =>'0', 115 =>'1', 116 =>'0', 117 =>'0', 118 =>'1', 119 =>'0', 
    120 =>'0', 121 =>'1', 122 =>'1', 123 =>'1', 124 =>'1', 125 =>'0', 126 =>'0', 127 =>'1', 128 =>'1', 129 =>'1', 
    130 =>'0', 131 =>'1', 132 =>'0', 133 =>'0', 134 =>'0', 135 =>'1', 136 =>'1', 137 =>'1', 138 =>'1', 139 =>'0', 
    140 =>'1', 141 =>'1', 142 =>'0', 143 =>'0', 144 =>'1', 145 =>'0', 146 =>'0'
  );

  constant vector2 : memory := 
  (
    0   =>'0', 1   =>'1', 2   =>'1', 3   =>'1', 4   =>'0', 5   =>'0', 6   =>'1', 7   =>'0', 8   =>'1', 9   =>'0', 
    10  =>'1', 11  =>'1', 12  =>'0', 13  =>'1', 14  =>'0', 15  =>'0', 16  =>'0', 17  =>'1', 18  =>'0', 19  =>'1', 
    20  =>'1', 21  =>'1', 22  =>'0', 23  =>'0', 24  =>'1', 25  =>'0', 26  =>'1', 27  =>'0', 28  =>'1', 29  =>'0', 
    30  =>'1', 31  =>'0', 32  =>'0', 33  =>'1', 34  =>'0', 35  =>'0', 36  =>'0', 37  =>'1', 38  =>'1', 39  =>'0', 
    40  =>'0', 41  =>'1', 42  =>'1', 43  =>'0', 44  =>'0', 45  =>'0', 46  =>'1', 47  =>'1', 48  =>'0', 49  =>'0',
    50  =>'1', 51  =>'1', 52  =>'0', 53  =>'1', 54  =>'1', 55  =>'0', 56  =>'1', 57  =>'1', 58  =>'1', 59  =>'0', 
    60  =>'0', 61  =>'1', 62  =>'0', 63  =>'0', 64  =>'1', 65  =>'0', 66  =>'0', 67  =>'1', 68  =>'0', 69  =>'0',
    70  =>'1', 71  =>'1', 72  =>'0', 73  =>'0', 74  =>'1', 75  =>'1', 76  =>'0', 77  =>'0', 78  =>'1', 79  =>'1', 
    80  =>'0', 81  =>'0', 82  =>'0', 83  =>'1', 84  =>'0', 85  =>'1', 86  =>'0', 87  =>'0', 88  =>'0', 89  =>'0', 
    90  =>'1', 91  =>'1', 92  =>'0', 93  =>'0', 94  =>'1', 95  =>'1', 96  =>'0', 97  =>'0', 98  =>'0', 99  =>'0',
    100 =>'1', 101 =>'0', 102 =>'1', 103 =>'1', 104 =>'1', 105 =>'1', 106 =>'0', 107 =>'0', 108 =>'0', 109 =>'1', 
    110 =>'1', 111 =>'0', 112 =>'0', 113 =>'1', 114 =>'0', 115 =>'1', 116 =>'0', 117 =>'1', 118 =>'1', 119 =>'0', 
    120 =>'1', 121 =>'1', 122 =>'1', 123 =>'1', 124 =>'1', 125 =>'0', 126 =>'1', 127 =>'1', 128 =>'0', 129 =>'0', 
    130 =>'0', 131 =>'0', 132 =>'0', 133 =>'1', 134 =>'0', 135 =>'1', 136 =>'0', 137 =>'1', 138 =>'0', 139 =>'0', 
    140 =>'0', 141 =>'0', 142 =>'0', 143 =>'1', 144 =>'1', 145 =>'0', 146 =>'0'
  );

  constant vector3 : memory := 
  (
    0   =>'0', 1   =>'1', 2   =>'1', 3   =>'0', 4   =>'1', 5   =>'1', 6   =>'0', 7   =>'0', 8   =>'1', 9   =>'0', 
    10  =>'1', 11  =>'1', 12  =>'1', 13  =>'1', 14  =>'0', 15  =>'1', 16  =>'0', 17  =>'1', 18  =>'1', 19  =>'1', 
    20  =>'0', 21  =>'1', 22  =>'1', 23  =>'1', 24  =>'1', 25  =>'0', 26  =>'1', 27  =>'0', 28  =>'1', 29  =>'0', 
    30  =>'1', 31  =>'1', 32  =>'0', 33  =>'1', 34  =>'0', 35  =>'1', 36  =>'0', 37  =>'1', 38  =>'1', 39  =>'0', 
    40  =>'0', 41  =>'0', 42  =>'1', 43  =>'0', 44  =>'1', 45  =>'0', 46  =>'1', 47  =>'1', 48  =>'0', 49  =>'0',
    50  =>'1', 51  =>'0', 52  =>'1', 53  =>'0', 54  =>'1', 55  =>'0', 56  =>'1', 57  =>'1', 58  =>'1', 59  =>'0', 
    60  =>'1', 61  =>'1', 62  =>'0', 63  =>'0', 64  =>'1', 65  =>'0', 66  =>'1', 67  =>'0', 68  =>'0', 69  =>'1',
    70  =>'1', 71  =>'0', 72  =>'1', 73  =>'1', 74  =>'0', 75  =>'1', 76  =>'1', 77  =>'1', 78  =>'0', 79  =>'0', 
    80  =>'1', 81  =>'0', 82  =>'0', 83  =>'1', 84  =>'1', 85  =>'0', 86  =>'1', 87  =>'0', 88  =>'1', 89  =>'1',
    90  =>'0', 91  =>'0', 92  =>'1', 93  =>'0', 94  =>'0', 95  =>'0', 96  =>'1', 97  =>'0', 98  =>'0', 99  =>'0',
    100 =>'1', 101 =>'0', 102 =>'1', 103 =>'1', 104 =>'1', 105 =>'1', 106 =>'0', 107 =>'0', 108 =>'0', 109 =>'1', 
    110 =>'0', 111 =>'0', 112 =>'1', 113 =>'0', 114 =>'0', 115 =>'1', 116 =>'0', 117 =>'1', 118 =>'1', 119 =>'0', 
    120 =>'1', 121 =>'1', 122 =>'1', 123 =>'1', 124 =>'1', 125 =>'0', 126 =>'1', 127 =>'1', 128 =>'0', 129 =>'0', 
    130 =>'0', 131 =>'0', 132 =>'0', 133 =>'1', 134 =>'0', 135 =>'1', 136 =>'0', 137 =>'1', 138 =>'0', 139 =>'0', 
    140 =>'0', 141 =>'1', 142 =>'0', 143 =>'0', 144 =>'1', 145 =>'0', 146 =>'0'
  );

  constant vector4 : memory := 
  (
    0   =>'0', 1   =>'0', 2   =>'1', 3   =>'0', 4   =>'1', 5   =>'0', 6   =>'0', 7   =>'0', 8   =>'0', 9   =>'0', 
    10  =>'1', 11  =>'0', 12  =>'1', 13  =>'1', 14  =>'0', 15  =>'1', 16  =>'0', 17  =>'1', 18  =>'1', 19  =>'0', 
    20  =>'0', 21  =>'1', 22  =>'1', 23  =>'1', 24  =>'1', 25  =>'0', 26  =>'1', 27  =>'1', 28  =>'1', 29  =>'0', 
    30  =>'1', 31  =>'0', 32  =>'0', 33  =>'1', 34  =>'0', 35  =>'1', 36  =>'1', 37  =>'1', 38  =>'1', 39  =>'1', 
    40  =>'0', 41  =>'0', 42  =>'1', 43  =>'0', 44  =>'1', 45  =>'0', 46  =>'1', 47  =>'1', 48  =>'0', 49  =>'0',
    50  =>'1', 51  =>'1', 52  =>'0', 53  =>'1', 54  =>'1', 55  =>'0', 56  =>'1', 57  =>'1', 58  =>'1', 59  =>'0', 
    60  =>'0', 61  =>'1', 62  =>'0', 63  =>'0', 64  =>'1', 65  =>'0', 66  =>'0', 67  =>'1', 68  =>'1', 69  =>'0',
    70  =>'0', 71  =>'0', 72  =>'1', 73  =>'1', 74  =>'0', 75  =>'1', 76  =>'1', 77  =>'1', 78  =>'0', 79  =>'0', 
    80  =>'1', 81  =>'1', 82  =>'1', 83  =>'0', 84  =>'0', 85  =>'1', 86  =>'0', 87  =>'0', 88  =>'1', 89  =>'1',
    90  =>'0', 91  =>'0', 92  =>'1', 93  =>'1', 94  =>'0', 95  =>'0', 96  =>'1', 97  =>'0', 98  =>'0', 99  =>'0',
    100 =>'1', 101 =>'0', 102 =>'1', 103 =>'1', 104 =>'1', 105 =>'1', 106 =>'1', 107 =>'0', 108 =>'0', 109 =>'1', 
    110 =>'0', 111 =>'0', 112 =>'1', 113 =>'0', 114 =>'1', 115 =>'1', 116 =>'1', 117 =>'0', 118 =>'1', 119 =>'0', 
    120 =>'0', 121 =>'1', 122 =>'1', 123 =>'0', 124 =>'1', 125 =>'0', 126 =>'1', 127 =>'1', 128 =>'1', 129 =>'0', 
    130 =>'1', 131 =>'0', 132 =>'0', 133 =>'1', 134 =>'0', 135 =>'1', 136 =>'1', 137 =>'1', 138 =>'0', 139 =>'0', 
    140 =>'0', 141 =>'1', 142 =>'1', 143 =>'0', 144 =>'1', 145 =>'0', 146 =>'0'
  );

  constant vector5 : memory := 
  (
    0   =>'0', 1   =>'1', 2   =>'1', 3   =>'0', 4   =>'1', 5   =>'1', 6   =>'0', 7   =>'0', 8   =>'1', 9   =>'0', 
    10  =>'1', 11  =>'0', 12  =>'1', 13  =>'1', 14  =>'0', 15  =>'1', 16  =>'0', 17  =>'1', 18  =>'1', 19  =>'1', 
    20  =>'0', 21  =>'1', 22  =>'1', 23  =>'1', 24  =>'1', 25  =>'0', 26  =>'1', 27  =>'0', 28  =>'1', 29  =>'0', 
    30  =>'1', 31  =>'1', 32  =>'0', 33  =>'1', 34  =>'0', 35  =>'1', 36  =>'0', 37  =>'1', 38  =>'1', 39  =>'0', 
    40  =>'0', 41  =>'0', 42  =>'1', 43  =>'0', 44  =>'1', 45  =>'0', 46  =>'1', 47  =>'1', 48  =>'0', 49  =>'0',
    50  =>'1', 51  =>'1', 52  =>'0', 53  =>'1', 54  =>'1', 55  =>'0', 56  =>'0', 57  =>'1', 58  =>'0', 59  =>'1', 
    60  =>'1', 61  =>'0', 62  =>'1', 63  =>'0', 64  =>'0', 65  =>'1', 66  =>'1', 67  =>'0', 68  =>'0', 69  =>'1', 
    70  =>'1', 71  =>'1', 72  =>'1', 73  =>'0', 74  =>'1', 75  =>'1', 76  =>'0', 77  =>'0', 78  =>'1', 79  =>'1', 
    80  =>'0', 81  =>'0', 82  =>'0', 83  =>'1', 84  =>'1', 85  =>'0', 86  =>'0', 87  =>'1', 88  =>'0', 89  =>'0',
    90  =>'1', 91  =>'1', 92  =>'0', 93  =>'0', 94  =>'1', 95  =>'0', 96  =>'0', 97  =>'0', 98  =>'0', 99  =>'1',
    100 =>'0', 101 =>'0', 102 =>'1', 103 =>'1', 104 =>'1', 105 =>'1', 106 =>'0', 107 =>'0', 108 =>'0', 109 =>'1', 
    110 =>'0', 111 =>'1', 112 =>'1', 113 =>'0', 114 =>'0', 115 =>'1', 116 =>'1', 117 =>'0', 118 =>'1', 119 =>'0', 
    120 =>'0', 121 =>'1', 122 =>'0', 123 =>'0', 124 =>'0', 125 =>'0', 126 =>'1', 127 =>'1', 128 =>'1', 129 =>'0', 
    130 =>'1', 131 =>'0', 132 =>'0', 133 =>'1', 134 =>'0', 135 =>'0', 136 =>'1', 137 =>'0', 138 =>'0', 139 =>'1', 
    140 =>'0', 141 =>'0', 142 =>'1', 143 =>'0', 144 =>'1', 145 =>'0', 146 =>'0'
  );

  constant vector6 : memory := 
  (
    0   =>'0', 1   =>'0', 2   =>'0', 3   =>'0', 4   =>'0', 5   =>'0', 6   =>'0', 7   =>'0', 8   =>'0', 9   =>'0', 
    10  =>'0', 11  =>'0', 12  =>'0', 13  =>'0', 14  =>'0', 15  =>'0', 16  =>'0', 17  =>'0', 18  =>'0', 19  =>'0', 
    20  =>'0', 21  =>'0', 22  =>'0', 23  =>'0', 24  =>'0', 25  =>'0', 26  =>'0', 27  =>'0', 28  =>'0', 29  =>'0', 
    30  =>'0', 31  =>'0', 32  =>'0', 33  =>'0', 34  =>'0', 35  =>'0', 36  =>'0', 37  =>'0', 38  =>'0', 39  =>'0', 
    40  =>'0', 41  =>'0', 42  =>'0', 43  =>'0', 44  =>'0', 45  =>'0', 46  =>'0', 47  =>'0', 48  =>'0', 49  =>'1', 
    50  =>'1', 51  =>'1', 52  =>'1', 53  =>'1', 54  =>'1', 55  =>'1', 56  =>'1', 57  =>'1', 58  =>'1', 59  =>'1', 
    60  =>'1', 61  =>'1', 62  =>'1', 63  =>'1', 64  =>'1', 65  =>'1', 66  =>'1', 67  =>'1', 68  =>'1', 69  =>'1',
    70  =>'1', 71  =>'1', 72  =>'1', 73  =>'1', 74  =>'1', 75  =>'1', 76  =>'1', 77  =>'1', 78  =>'1', 79  =>'1', 
    80  =>'1', 81  =>'1', 82  =>'1', 83  =>'1', 84  =>'1', 85  =>'1', 86  =>'1', 87  =>'1', 88  =>'1', 89  =>'1',
    90  =>'1', 91  =>'1', 92  =>'1', 93  =>'1', 94  =>'1', 95  =>'1', 96  =>'1', 97  =>'0', 98  =>'0', 99  =>'0', 
    100 =>'0', 101 =>'0', 102 =>'0', 103 =>'0', 104 =>'0', 105 =>'0', 106 =>'0', 107 =>'0', 108 =>'0', 109 =>'0', 
    110 =>'0', 111 =>'0', 112 =>'0', 113 =>'0', 114 =>'0', 115 =>'0', 116 =>'0', 117 =>'0', 118 =>'0', 119 =>'0', 
    120 =>'0', 121 =>'0', 122 =>'0', 123 =>'0', 124 =>'0', 125 =>'0', 126 =>'0', 127 =>'0', 128 =>'0', 129 =>'0', 
    130 =>'0', 131 =>'0', 132 =>'0', 133 =>'0', 134 =>'0', 135 =>'0', 136 =>'0', 137 =>'0', 138 =>'0', 139 =>'0', 
    140 =>'0', 141 =>'0', 142 =>'0', 143 =>'0', 144 =>'0', 145 =>'0', 146 =>'0'
  );

begin 
   
  process(clk) is
  begin 
    if rising_edge(clk) then 
      data1 <= vector1(to_integer(unsigned(address)));
      data2 <= vector2(to_integer(unsigned(address)));
      data3 <= vector3(to_integer(unsigned(address)));
      data4 <= vector4(to_integer(unsigned(address)));
      data5 <= vector5(to_integer(unsigned(address)));
      data6 <= vector6(to_integer(unsigned(address)));
    end if;
  end process;
  
end architecture;
